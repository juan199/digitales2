
module transmitter(
	input wire       TXCLK,
	input wire       INTERCLK,
	input wire       TRANSCLK,
	input wire [7:0] TXDATA,
	input wire       TXDATAK,
	input wire       TXCOMP,
	input wire       DATALOOPB,
	input wire       RXLOOPB,
	input wire       TXIDEL,
	input wire       TXDET,
	output wire      RXDET_O,
	output wire      TX_P,
	output wire      TX_N	
);


endmodule
