module bancodepruebas;
	codificador conducta(S1,S2,S3,S4,E1,E2,E3,E4);
	probador pruebas(S1,S2,S3,S4,S1e,S2e,S3e,S4e,E1,E2,E3,E4);
	cod_str estructural(S1e,S2e,S3e,S4e,E1,E2,E3,E4);
endmodule